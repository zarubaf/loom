// SPDX-License-Identifier: Apache-2.0
// Loom Scan Chain Controller
//
// Controls scan chain capture (shift out state) and restore (shift in state).
// With free-running clock + FF enable override (loom_en | loom_scan_enable),
// the scan controller simply asserts scan_enable and shifts one bit per cycle.
//
// Register Map (offset from base):
//   0x00 SCAN_STATUS    R    [0]=busy, [1]=done, [7:4]=error_code
//   0x04 SCAN_CONTROL   W    Command: 1=capture, 2=restore
//   0x08 SCAN_LENGTH    R    Chain length in bits (from parameter)
//   0x0C reserved
//   0x10 SCAN_DATA[0]   RW   First 32 bits of scan data (LSBs)
//   0x14 SCAN_DATA[1]   RW   Next 32 bits
//   ...
//
// Scan data is stored LSB-first: DATA[0][0] is the first bit shifted out/in.
// Maximum supported chain length is 32 * N_DATA_WORDS bits.

module loom_scan_ctrl #(
    parameter int unsigned CHAIN_LENGTH  = 64,   // Total scan chain bits
    parameter int unsigned N_DATA_WORDS  = (CHAIN_LENGTH + 31) / 32  // Data buffer size
)(
    input  logic        clk_i,
    input  logic        rst_ni,

    // AXI-Lite Slave interface
    input  logic [11:0] axil_araddr_i,
    input  logic        axil_arvalid_i,
    output logic        axil_arready_o,
    output logic [31:0] axil_rdata_o,
    output logic [1:0]  axil_rresp_o,
    output logic        axil_rvalid_o,
    input  logic        axil_rready_i,

    input  logic [11:0] axil_awaddr_i,
    input  logic        axil_awvalid_i,
    output logic        axil_awready_o,
    input  logic [31:0] axil_wdata_i,
    input  logic        axil_wvalid_i,
    output logic        axil_wready_o,
    output logic [1:0]  axil_bresp_o,
    output logic        axil_bvalid_o,
    input  logic        axil_bready_i,

    // Scan chain interface (directly to DUT)
    output logic        scan_enable_o,    // Scan mode enable (to loom_scan_enable)
    output logic        scan_in_o,        // Serial data in (to loom_scan_in)
    input  logic        scan_out_i,       // Serial data out (from loom_scan_out)

    // Status output
    output logic        scan_busy_o       // Scan operation in progress
);

    // =========================================================================
    // State Machine
    // =========================================================================

    typedef enum logic [2:0] {
        StIdle     = 3'd0,
        StCapture  = 3'd1,  // Shifting data out of scan chain
        StRestore  = 3'd2,  // Shifting data into scan chain
        StDone     = 3'd3
    } state_e;

    // Command codes
    localparam logic [7:0] CMD_CAPTURE = 8'h01;
    localparam logic [7:0] CMD_RESTORE = 8'h02;

    // Widths for bit position / word index — avoid degenerate zero-width signals
    localparam int unsigned SHIFT_CNT_W = $clog2(CHAIN_LENGTH + 1);
    localparam int unsigned BIT_POS_W   = (CHAIN_LENGTH > 1) ? $clog2(CHAIN_LENGTH) : 1;

    state_e state_q;
    logic [SHIFT_CNT_W-1:0] shift_count_q;  // Bits remaining to shift
    logic [31:0] scan_data_q [N_DATA_WORDS]; // Scan data buffer
    logic        done_q;                     // Operation completed
    logic [3:0]  error_code_q;

    // =========================================================================
    // Scan Shift Logic
    // =========================================================================

    // Current bit position in the data buffer.
    // shift_count_q counts down from CHAIN_LENGTH.  We number buffer positions
    // so that position 0 corresponds to the LAST bit shifted out (= the bit
    // closest to scan_in, i.e. the first FF's LSB).  This matches the offset
    // numbering in the scan_map generated by scan_insert.
    logic [BIT_POS_W-1:0] bit_pos;
    assign bit_pos = BIT_POS_W'(shift_count_q) - BIT_POS_W'(1);

    // Which word and bit within that word
    logic [4:0] bit_in_word;
    assign bit_in_word = bit_pos[4:0];

    // Word index: bit_pos / 32.  For single-word chains, always 0.
    logic [$clog2(N_DATA_WORDS > 1 ? N_DATA_WORDS : 2)-1:0] word_idx;
    generate
        if (N_DATA_WORDS > 1)
            assign word_idx = bit_pos[BIT_POS_W-1:5];
        else
            assign word_idx = '0;
    endgenerate

    // Scan input data:
    //   Capture: closed-loop — feed scan_out back to scan_in so the chain
    //           contents are preserved after a full capture (non-destructive).
    //   Restore: feed from the data buffer to overwrite chain contents.
    assign scan_in_o = (state_q == StCapture)  ? scan_out_i :
                       (state_q == StRestore && shift_count_q > 0) ?
                       scan_data_q[word_idx][bit_in_word] : 1'b0;

    // Scan enable: active during capture or restore, but only while shifts remain.
    // Without the shift_count_q guard, an extra shift occurs on the cycle where
    // shift_count_q == 0 (state_q hasn't transitioned to StDone yet).
    assign scan_enable_o = (state_q == StCapture || state_q == StRestore)
                           && (shift_count_q != '0);

    // Busy output
    assign scan_busy_o = (state_q != StIdle && state_q != StDone);

    // =========================================================================
    // AXI-Lite Write Handshake
    // =========================================================================

    logic        wr_addr_valid_q, wr_data_valid_q;
    logic [11:0] wr_addr_q;
    logic [31:0] wr_data_q;

    // Write-effect decode (combinational) — consumed by main FSM
    logic       wr_fire;       // write handshake fires this cycle
    logic       wr_cmd_capture;
    logic       wr_cmd_restore;
    logic       wr_clear_done;
    logic       wr_data_en;
    logic [9:0] wr_data_word_addr;

    assign wr_fire = wr_addr_valid_q && wr_data_valid_q && !axil_bvalid_o;

    always_comb begin
        wr_cmd_capture   = 1'b0;
        wr_cmd_restore   = 1'b0;
        wr_clear_done    = 1'b0;
        wr_data_en       = 1'b0;
        wr_data_word_addr = '0;

        if (wr_fire) begin
            case (wr_addr_q[11:2])
                10'h000: begin  // SCAN_STATUS — write-to-clear done
                    wr_clear_done = wr_data_q[1];
                end
                10'h001: begin  // SCAN_CONTROL
                    case (wr_data_q[7:0])
                        CMD_CAPTURE: wr_cmd_capture = 1'b1;
                        CMD_RESTORE: wr_cmd_restore = 1'b1;
                        default: ;
                    endcase
                end
                default: begin
                    // SCAN_DATA registers (offset 0x10 = word address 4)
                    if (wr_addr_q[11:2] >= 10'h004 &&
                        wr_addr_q[11:2] < 10'h004 + N_DATA_WORDS[9:0]) begin
                        wr_data_en       = 1'b1;
                        wr_data_word_addr = wr_addr_q[11:2] - 10'h004;
                    end
                end
            endcase
        end
    end

    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            wr_addr_valid_q <= 1'b0;
            wr_data_valid_q <= 1'b0;
            wr_addr_q       <= 12'd0;
            wr_data_q       <= 32'd0;
            axil_awready_o  <= 1'b0;
            axil_wready_o   <= 1'b0;
            axil_bvalid_o   <= 1'b0;
            axil_bresp_o    <= 2'b00;
        end else begin
            axil_awready_o <= 1'b1;
            axil_wready_o  <= 1'b1;

            if (axil_awvalid_i && axil_awready_o) begin
                wr_addr_q       <= axil_awaddr_i;
                wr_addr_valid_q <= 1'b1;
            end

            if (axil_wvalid_i && axil_wready_o) begin
                wr_data_q       <= axil_wdata_i;
                wr_data_valid_q <= 1'b1;
            end

            if (wr_fire) begin
                wr_addr_valid_q <= 1'b0;
                wr_data_valid_q <= 1'b0;
                axil_bvalid_o   <= 1'b1;
                axil_bresp_o    <= 2'b00;
            end

            if (axil_bvalid_o && axil_bready_i) begin
                axil_bvalid_o <= 1'b0;
            end
        end
    end

    // =========================================================================
    // Main FSM — single always_ff block (no multi-driven signals)
    // =========================================================================

    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            state_q       <= StIdle;
            shift_count_q <= '0;
            done_q        <= 1'b0;
            error_code_q  <= 4'd0;
            for (int i = 0; i < int'(N_DATA_WORDS); i++) begin
                scan_data_q[i] <= 32'd0;
            end
        end else begin
            case (state_q)
                StIdle: begin
                    // Write effects while idle
                    if (wr_cmd_capture) begin
                        state_q       <= StCapture;
                        shift_count_q <= SHIFT_CNT_W'(CHAIN_LENGTH);
                        done_q        <= 1'b0;
                        error_code_q  <= 4'd0;
                    end else if (wr_cmd_restore) begin
                        state_q       <= StRestore;
                        shift_count_q <= SHIFT_CNT_W'(CHAIN_LENGTH);
                        done_q        <= 1'b0;
                        error_code_q  <= 4'd0;
                    end
                    if (wr_clear_done) begin
                        done_q <= 1'b0;
                    end
                    if (wr_data_en) begin
                        scan_data_q[wr_data_word_addr] <= wr_data_q;
                    end
                end

                StCapture: begin
                    if (shift_count_q > 0) begin
                        scan_data_q[word_idx][bit_in_word] <= scan_out_i;
                        shift_count_q <= shift_count_q - 1;
                    end else begin
                        state_q <= StDone;
                    end
                end

                StRestore: begin
                    if (shift_count_q > 0) begin
                        shift_count_q <= shift_count_q - 1;
                    end else begin
                        state_q <= StDone;
                    end
                end

                StDone: begin
                    done_q <= 1'b1;
                    // Write effects while done
                    if (wr_clear_done) begin
                        done_q  <= 1'b0;
                        state_q <= StIdle;
                    end
                    if (wr_data_en) begin
                        scan_data_q[wr_data_word_addr] <= wr_data_q;
                    end
                end

                default: state_q <= StIdle;
            endcase
        end
    end

    // =========================================================================
    // AXI-Lite Read Interface
    // =========================================================================

    logic [11:0] rd_addr_q;
    logic        rd_pending_q;

    always_ff @(posedge clk_i or negedge rst_ni) begin
        if (!rst_ni) begin
            rd_pending_q   <= 1'b0;
            rd_addr_q      <= 12'd0;
            axil_arready_o <= 1'b0;
            axil_rvalid_o  <= 1'b0;
            axil_rdata_o   <= 32'd0;
            axil_rresp_o   <= 2'b00;
        end else begin
            axil_arready_o <= 1'b1;

            if (axil_arvalid_i && axil_arready_o) begin
                rd_addr_q    <= axil_araddr_i;
                rd_pending_q <= 1'b1;
            end

            if (rd_pending_q && !axil_rvalid_o) begin
                axil_rvalid_o <= 1'b1;
                axil_rresp_o  <= 2'b00;

                case (rd_addr_q[11:2])
                    10'h000: axil_rdata_o <= {24'd0, error_code_q, 2'd0, done_q, scan_busy_o};  // SCAN_STATUS
                    10'h002: axil_rdata_o <= CHAIN_LENGTH;  // SCAN_LENGTH
                    default: begin
                        // SCAN_DATA registers start at offset 0x10 (word address 4)
                        if (rd_addr_q[11:2] >= 10'h004 &&
                            rd_addr_q[11:2] < 10'h004 + N_DATA_WORDS[9:0]) begin
                            axil_rdata_o <= scan_data_q[rd_addr_q[11:2] - 10'h004];
                        end else begin
                            axil_rdata_o <= 32'hDEAD_BEEF;
                        end
                    end
                endcase

                rd_pending_q <= 1'b0;
            end

            if (axil_rvalid_o && axil_rready_i) begin
                axil_rvalid_o <= 1'b0;
            end
        end
    end

endmodule
