// SPDX-License-Identifier: Apache-2.0
// tb_emu_top.sv - End-to-end testbench for emulation wrapper
//
// This testbench demonstrates the full emu_top flow:
// 1. emu_top wrapper with clock gating
// 2. loom_host_stub handling DPI calls
// 3. Design execution with automatic clock gate/release

`timescale 1ns/1ps

module tb_emu_top;

    // Clock and reset
    logic clk;
    logic rst;

    // DUT interface signals
    logic [31:0] a, b;
    logic start;
    logic [31:0] result;
    logic done;

    // DPI interface (directly from wrapper)
    logic        dpi_valid;
    logic        dpi_ack;
    logic [7:0]  dpi_func_id;
    logic [63:0] dpi_args;
    logic [31:0] dpi_result;

    // Scan interface
    logic scan_enable;
    logic scan_in;
    logic scan_out;

    // Clock generation (100 MHz)
    initial clk = 0;
    always #5 clk = ~clk;

    // Instantiate the emu_top wrapper (generated by Yosys)
    emu_top_dpi_example u_emu_top (
        .clk              (clk),
        .rst              (rst),
        .a                (a),
        .b                (b),
        .start            (start),
        .result           (result),
        .done             (done),
        .loom_dpi_valid   (dpi_valid),
        .loom_dpi_ack     (dpi_ack),
        .loom_dpi_func_id (dpi_func_id),
        .loom_dpi_args    (dpi_args),
        .loom_dpi_result  (dpi_result),
        .loom_scan_enable (scan_enable),
        .loom_scan_in     (scan_in),
        .loom_scan_out    (scan_out)
    );

    // Instantiate host stub to handle DPI calls
    loom_host_stub #(
        .FUNC_ID_WIDTH (8),
        .MAX_ARG_WIDTH (64),
        .MAX_RET_WIDTH (32),
        .HOST_LATENCY  (0)  // 0 cycle latency for faster simulation
    ) u_host_stub (
        .clk        (clk),
        .rst        (rst),
        .dpi_valid  (dpi_valid),
        .dpi_func_id(dpi_func_id),
        .dpi_args   (dpi_args),
        .dpi_result (dpi_result),
        .dpi_ack    (dpi_ack)
    );

    // Test sequence
    initial begin
        $dumpfile("tb_emu_top.vcd");
        $dumpvars(0, tb_emu_top);

        // Initialize
        rst = 1;
        a = 0;
        b = 0;
        start = 0;
        scan_enable = 0;
        scan_in = 0;

        // Reset sequence
        repeat (10) @(posedge clk);
        rst = 0;
        repeat (5) @(posedge clk);

        $display("\n=== Test 1: DPI addition (10 + 20) ===");
        a = 32'd10;
        b = 32'd20;
        start = 1;
        @(posedge clk);
        start = 0;

        // Wait for done (DPI call will gate clock, host stub will respond)
        wait(done);
        @(posedge clk);

        if (result == 32'd30) begin
            $display("PASS: result = %0d (expected 30)", result);
        end else begin
            $display("FAIL: result = %0d (expected 30)", result);
        end

        repeat (10) @(posedge clk);

        $display("\n=== Test 2: DPI addition (100 + 200) ===");
        a = 32'd100;
        b = 32'd200;
        start = 1;
        @(posedge clk);
        start = 0;

        wait(done);
        @(posedge clk);

        if (result == 32'd300) begin
            $display("PASS: result = %0d (expected 300)", result);
        end else begin
            $display("FAIL: result = %0d (expected 300)", result);
        end

        repeat (10) @(posedge clk);

        $display("\n=== All tests complete ===");
        $finish;
    end

    // Timeout watchdog
    initial begin
        #50000;
        $display("ERROR: Timeout - simulation did not complete");
        $finish;
    end

    // Monitor clock gating
    always @(posedge clk) begin
        if (!rst && dpi_valid && !dpi_ack) begin
            $display("[%0t] Clock GATED - DPI call pending: func_id=%0d, args=%h", $time, dpi_func_id, dpi_args);
        end
    end

    always @(posedge dpi_ack) begin
        if (!rst) begin
            $display("[%0t] Clock RELEASED - Host ACK, result: %0d", $time, dpi_result);
        end
    end

endmodule
